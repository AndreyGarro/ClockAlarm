// clock.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module clock (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] cpu_data_master_readdata;                          // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                       // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                       // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [13:0] cpu_data_master_address;                           // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                        // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                              // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                             // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                         // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                   // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [13:0] cpu_instruction_master_address;                    // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                       // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;    // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest; // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess; // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;     // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;        // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;  // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;       // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;   // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;               // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                 // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_s1_address;                  // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;               // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                    // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                    // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_reg_bu_s1_chipselect;            // mm_interconnect_0:REG_Bu_s1_chipselect -> REG_Bu:chipselect
	wire  [31:0] mm_interconnect_0_reg_bu_s1_readdata;              // REG_Bu:readdata -> mm_interconnect_0:REG_Bu_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_bu_s1_address;               // mm_interconnect_0:REG_Bu_s1_address -> REG_Bu:address
	wire         mm_interconnect_0_reg_bu_s1_write;                 // mm_interconnect_0:REG_Bu_s1_write -> REG_Bu:write_n
	wire  [31:0] mm_interconnect_0_reg_bu_s1_writedata;             // mm_interconnect_0:REG_Bu_s1_writedata -> REG_Bu:writedata
	wire         mm_interconnect_0_reg_bd_s1_chipselect;            // mm_interconnect_0:REG_Bd_s1_chipselect -> REG_Bd:chipselect
	wire  [31:0] mm_interconnect_0_reg_bd_s1_readdata;              // REG_Bd:readdata -> mm_interconnect_0:REG_Bd_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_bd_s1_address;               // mm_interconnect_0:REG_Bd_s1_address -> REG_Bd:address
	wire         mm_interconnect_0_reg_bd_s1_write;                 // mm_interconnect_0:REG_Bd_s1_write -> REG_Bd:write_n
	wire  [31:0] mm_interconnect_0_reg_bd_s1_writedata;             // mm_interconnect_0:REG_Bd_s1_writedata -> REG_Bd:writedata
	wire         mm_interconnect_0_reg_bn_s1_chipselect;            // mm_interconnect_0:REG_Bn_s1_chipselect -> REG_Bn:chipselect
	wire  [31:0] mm_interconnect_0_reg_bn_s1_readdata;              // REG_Bn:readdata -> mm_interconnect_0:REG_Bn_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_bn_s1_address;               // mm_interconnect_0:REG_Bn_s1_address -> REG_Bn:address
	wire         mm_interconnect_0_reg_bn_s1_write;                 // mm_interconnect_0:REG_Bn_s1_write -> REG_Bn:write_n
	wire  [31:0] mm_interconnect_0_reg_bn_s1_writedata;             // mm_interconnect_0:REG_Bn_s1_writedata -> REG_Bn:writedata
	wire         mm_interconnect_0_reg_bs_s1_chipselect;            // mm_interconnect_0:REG_Bs_s1_chipselect -> REG_Bs:chipselect
	wire  [31:0] mm_interconnect_0_reg_bs_s1_readdata;              // REG_Bs:readdata -> mm_interconnect_0:REG_Bs_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_bs_s1_address;               // mm_interconnect_0:REG_Bs_s1_address -> REG_Bs:address
	wire         mm_interconnect_0_reg_bs_s1_write;                 // mm_interconnect_0:REG_Bs_s1_write -> REG_Bs:write_n
	wire  [31:0] mm_interconnect_0_reg_bs_s1_writedata;             // mm_interconnect_0:REG_Bs_s1_writedata -> REG_Bs:writedata
	wire         mm_interconnect_0_reg_h1_s1_chipselect;            // mm_interconnect_0:REG_H1_s1_chipselect -> REG_H1:chipselect
	wire  [31:0] mm_interconnect_0_reg_h1_s1_readdata;              // REG_H1:readdata -> mm_interconnect_0:REG_H1_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_h1_s1_address;               // mm_interconnect_0:REG_H1_s1_address -> REG_H1:address
	wire         mm_interconnect_0_reg_h1_s1_write;                 // mm_interconnect_0:REG_H1_s1_write -> REG_H1:write_n
	wire  [31:0] mm_interconnect_0_reg_h1_s1_writedata;             // mm_interconnect_0:REG_H1_s1_writedata -> REG_H1:writedata
	wire         mm_interconnect_0_reg_h2_s1_chipselect;            // mm_interconnect_0:REG_H2_s1_chipselect -> REG_H2:chipselect
	wire  [31:0] mm_interconnect_0_reg_h2_s1_readdata;              // REG_H2:readdata -> mm_interconnect_0:REG_H2_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_h2_s1_address;               // mm_interconnect_0:REG_H2_s1_address -> REG_H2:address
	wire         mm_interconnect_0_reg_h2_s1_write;                 // mm_interconnect_0:REG_H2_s1_write -> REG_H2:write_n
	wire  [31:0] mm_interconnect_0_reg_h2_s1_writedata;             // mm_interconnect_0:REG_H2_s1_writedata -> REG_H2:writedata
	wire         mm_interconnect_0_reg_m1_s1_chipselect;            // mm_interconnect_0:REG_M1_s1_chipselect -> REG_M1:chipselect
	wire  [31:0] mm_interconnect_0_reg_m1_s1_readdata;              // REG_M1:readdata -> mm_interconnect_0:REG_M1_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_m1_s1_address;               // mm_interconnect_0:REG_M1_s1_address -> REG_M1:address
	wire         mm_interconnect_0_reg_m1_s1_write;                 // mm_interconnect_0:REG_M1_s1_write -> REG_M1:write_n
	wire  [31:0] mm_interconnect_0_reg_m1_s1_writedata;             // mm_interconnect_0:REG_M1_s1_writedata -> REG_M1:writedata
	wire         mm_interconnect_0_reg_m2_s1_chipselect;            // mm_interconnect_0:REG_M2_s1_chipselect -> REG_M2:chipselect
	wire  [31:0] mm_interconnect_0_reg_m2_s1_readdata;              // REG_M2:readdata -> mm_interconnect_0:REG_M2_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_m2_s1_address;               // mm_interconnect_0:REG_M2_s1_address -> REG_M2:address
	wire         mm_interconnect_0_reg_m2_s1_write;                 // mm_interconnect_0:REG_M2_s1_write -> REG_M2:write_n
	wire  [31:0] mm_interconnect_0_reg_m2_s1_writedata;             // mm_interconnect_0:REG_M2_s1_writedata -> REG_M2:writedata
	wire         mm_interconnect_0_reg_s1_s1_chipselect;            // mm_interconnect_0:REG_S1_s1_chipselect -> REG_S1:chipselect
	wire  [31:0] mm_interconnect_0_reg_s1_s1_readdata;              // REG_S1:readdata -> mm_interconnect_0:REG_S1_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_s1_s1_address;               // mm_interconnect_0:REG_S1_s1_address -> REG_S1:address
	wire         mm_interconnect_0_reg_s1_s1_write;                 // mm_interconnect_0:REG_S1_s1_write -> REG_S1:write_n
	wire  [31:0] mm_interconnect_0_reg_s1_s1_writedata;             // mm_interconnect_0:REG_S1_s1_writedata -> REG_S1:writedata
	wire         mm_interconnect_0_reg_s2_s1_chipselect;            // mm_interconnect_0:REG_S2_s1_chipselect -> REG_S2:chipselect
	wire  [31:0] mm_interconnect_0_reg_s2_s1_readdata;              // REG_S2:readdata -> mm_interconnect_0:REG_S2_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_s2_s1_address;               // mm_interconnect_0:REG_S2_s1_address -> REG_S2:address
	wire         mm_interconnect_0_reg_s2_s1_write;                 // mm_interconnect_0:REG_S2_s1_write -> REG_S2:write_n
	wire  [31:0] mm_interconnect_0_reg_s2_s1_writedata;             // mm_interconnect_0:REG_S2_s1_writedata -> REG_S2:writedata
	wire         mm_interconnect_0_reg_led_s1_chipselect;           // mm_interconnect_0:REG_LED_s1_chipselect -> REG_LED:chipselect
	wire  [31:0] mm_interconnect_0_reg_led_s1_readdata;             // REG_LED:readdata -> mm_interconnect_0:REG_LED_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_led_s1_address;              // mm_interconnect_0:REG_LED_s1_address -> REG_LED:address
	wire         mm_interconnect_0_reg_led_s1_write;                // mm_interconnect_0:REG_LED_s1_write -> REG_LED:write_n
	wire  [31:0] mm_interconnect_0_reg_led_s1_writedata;            // mm_interconnect_0:REG_LED_s1_writedata -> REG_LED:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;              // mm_interconnect_0:UART_s1_chipselect -> UART:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                // UART:readdata -> mm_interconnect_0:UART_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                 // mm_interconnect_0:UART_s1_address -> UART:address
	wire         mm_interconnect_0_uart_s1_read;                    // mm_interconnect_0:UART_s1_read -> UART:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;           // mm_interconnect_0:UART_s1_begintransfer -> UART:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                   // mm_interconnect_0:UART_s1_write -> UART:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;               // mm_interconnect_0:UART_s1_writedata -> UART:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;             // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;               // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                  // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;              // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         irq_mapper_receiver0_irq;                          // UART:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                          // REG_Bu:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                          // REG_Bd:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                          // REG_Bn:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                          // REG_Bs:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                          // TIMER:irq -> irq_mapper:receiver5_irq
	wire  [31:0] cpu_irq_irq;                                       // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                    // rst_controller:reset_out -> [CPU:reset_n, RAM:reset, REG_Bd:reset_n, REG_Bn:reset_n, REG_Bs:reset_n, REG_Bu:reset_n, REG_H1:reset_n, REG_H2:reset_n, REG_LED:reset_n, REG_M1:reset_n, REG_M2:reset_n, REG_S1:reset_n, REG_S2:reset_n, TIMER:reset_n, UART:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                // rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	clock_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	clock_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	clock_REG_Bd reg_bd (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_bd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_bd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_bd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_bd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_bd_s1_readdata),   //                    .readdata
		.in_port    (),                                       // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                //                 irq.irq
	);

	clock_REG_Bd reg_bn (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_bn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_bn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_bn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_bn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_bn_s1_readdata),   //                    .readdata
		.in_port    (),                                       // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                //                 irq.irq
	);

	clock_REG_Bd reg_bs (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_bs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_bs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_bs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_bs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_bs_s1_readdata),   //                    .readdata
		.in_port    (),                                       // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                //                 irq.irq
	);

	clock_REG_Bd reg_bu (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_bu_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_bu_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_bu_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_bu_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_bu_s1_readdata),   //                    .readdata
		.in_port    (),                                       // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                //                 irq.irq
	);

	clock_REG_H1 reg_h1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_h1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_h1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_h1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_h1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_h1_s1_readdata),   //                    .readdata
		.out_port   ()                                        // external_connection.export
	);

	clock_REG_H1 reg_h2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_h2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_h2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_h2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_h2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_h2_s1_readdata),   //                    .readdata
		.out_port   ()                                        // external_connection.export
	);

	clock_REG_H1 reg_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_reg_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_led_s1_readdata),   //                    .readdata
		.out_port   ()                                         // external_connection.export
	);

	clock_REG_H1 reg_m1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_m1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_m1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_m1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_m1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_m1_s1_readdata),   //                    .readdata
		.out_port   ()                                        // external_connection.export
	);

	clock_REG_H1 reg_m2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_m2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_m2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_m2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_m2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_m2_s1_readdata),   //                    .readdata
		.out_port   ()                                        // external_connection.export
	);

	clock_REG_H1 reg_s1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_s1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_s1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_s1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_s1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_s1_s1_readdata),   //                    .readdata
		.out_port   ()                                        // external_connection.export
	);

	clock_REG_H1 reg_s2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_s2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_s2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_s2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_s2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_s2_s1_readdata),   //                    .readdata
		.out_port   ()                                        // external_connection.export
	);

	clock_TIMER timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)               //   irq.irq
	);

	clock_UART uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (),                                        // external_connection.export
		.txd           (),                                        //                    .export
		.irq           (irq_mapper_receiver0_irq)                 //                 irq.irq
	);

	clock_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                           (clk_clk),                                           //                         CLK_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // CPU_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address               (cpu_data_master_address),                           //                 CPU_data_master.address
		.CPU_data_master_waitrequest           (cpu_data_master_waitrequest),                       //                                .waitrequest
		.CPU_data_master_byteenable            (cpu_data_master_byteenable),                        //                                .byteenable
		.CPU_data_master_read                  (cpu_data_master_read),                              //                                .read
		.CPU_data_master_readdata              (cpu_data_master_readdata),                          //                                .readdata
		.CPU_data_master_write                 (cpu_data_master_write),                             //                                .write
		.CPU_data_master_writedata             (cpu_data_master_writedata),                         //                                .writedata
		.CPU_data_master_debugaccess           (cpu_data_master_debugaccess),                       //                                .debugaccess
		.CPU_instruction_master_address        (cpu_instruction_master_address),                    //          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                //                                .waitrequest
		.CPU_instruction_master_read           (cpu_instruction_master_read),                       //                                .read
		.CPU_instruction_master_readdata       (cpu_instruction_master_readdata),                   //                                .readdata
		.CPU_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),     //             CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),       //                                .write
		.CPU_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),        //                                .read
		.CPU_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                                .readdata
		.CPU_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                                .writedata
		.CPU_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                                .byteenable
		.CPU_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                                .waitrequest
		.CPU_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                                .debugaccess
		.RAM_s1_address                        (mm_interconnect_0_ram_s1_address),                  //                          RAM_s1.address
		.RAM_s1_write                          (mm_interconnect_0_ram_s1_write),                    //                                .write
		.RAM_s1_readdata                       (mm_interconnect_0_ram_s1_readdata),                 //                                .readdata
		.RAM_s1_writedata                      (mm_interconnect_0_ram_s1_writedata),                //                                .writedata
		.RAM_s1_byteenable                     (mm_interconnect_0_ram_s1_byteenable),               //                                .byteenable
		.RAM_s1_chipselect                     (mm_interconnect_0_ram_s1_chipselect),               //                                .chipselect
		.RAM_s1_clken                          (mm_interconnect_0_ram_s1_clken),                    //                                .clken
		.REG_Bd_s1_address                     (mm_interconnect_0_reg_bd_s1_address),               //                       REG_Bd_s1.address
		.REG_Bd_s1_write                       (mm_interconnect_0_reg_bd_s1_write),                 //                                .write
		.REG_Bd_s1_readdata                    (mm_interconnect_0_reg_bd_s1_readdata),              //                                .readdata
		.REG_Bd_s1_writedata                   (mm_interconnect_0_reg_bd_s1_writedata),             //                                .writedata
		.REG_Bd_s1_chipselect                  (mm_interconnect_0_reg_bd_s1_chipselect),            //                                .chipselect
		.REG_Bn_s1_address                     (mm_interconnect_0_reg_bn_s1_address),               //                       REG_Bn_s1.address
		.REG_Bn_s1_write                       (mm_interconnect_0_reg_bn_s1_write),                 //                                .write
		.REG_Bn_s1_readdata                    (mm_interconnect_0_reg_bn_s1_readdata),              //                                .readdata
		.REG_Bn_s1_writedata                   (mm_interconnect_0_reg_bn_s1_writedata),             //                                .writedata
		.REG_Bn_s1_chipselect                  (mm_interconnect_0_reg_bn_s1_chipselect),            //                                .chipselect
		.REG_Bs_s1_address                     (mm_interconnect_0_reg_bs_s1_address),               //                       REG_Bs_s1.address
		.REG_Bs_s1_write                       (mm_interconnect_0_reg_bs_s1_write),                 //                                .write
		.REG_Bs_s1_readdata                    (mm_interconnect_0_reg_bs_s1_readdata),              //                                .readdata
		.REG_Bs_s1_writedata                   (mm_interconnect_0_reg_bs_s1_writedata),             //                                .writedata
		.REG_Bs_s1_chipselect                  (mm_interconnect_0_reg_bs_s1_chipselect),            //                                .chipselect
		.REG_Bu_s1_address                     (mm_interconnect_0_reg_bu_s1_address),               //                       REG_Bu_s1.address
		.REG_Bu_s1_write                       (mm_interconnect_0_reg_bu_s1_write),                 //                                .write
		.REG_Bu_s1_readdata                    (mm_interconnect_0_reg_bu_s1_readdata),              //                                .readdata
		.REG_Bu_s1_writedata                   (mm_interconnect_0_reg_bu_s1_writedata),             //                                .writedata
		.REG_Bu_s1_chipselect                  (mm_interconnect_0_reg_bu_s1_chipselect),            //                                .chipselect
		.REG_H1_s1_address                     (mm_interconnect_0_reg_h1_s1_address),               //                       REG_H1_s1.address
		.REG_H1_s1_write                       (mm_interconnect_0_reg_h1_s1_write),                 //                                .write
		.REG_H1_s1_readdata                    (mm_interconnect_0_reg_h1_s1_readdata),              //                                .readdata
		.REG_H1_s1_writedata                   (mm_interconnect_0_reg_h1_s1_writedata),             //                                .writedata
		.REG_H1_s1_chipselect                  (mm_interconnect_0_reg_h1_s1_chipselect),            //                                .chipselect
		.REG_H2_s1_address                     (mm_interconnect_0_reg_h2_s1_address),               //                       REG_H2_s1.address
		.REG_H2_s1_write                       (mm_interconnect_0_reg_h2_s1_write),                 //                                .write
		.REG_H2_s1_readdata                    (mm_interconnect_0_reg_h2_s1_readdata),              //                                .readdata
		.REG_H2_s1_writedata                   (mm_interconnect_0_reg_h2_s1_writedata),             //                                .writedata
		.REG_H2_s1_chipselect                  (mm_interconnect_0_reg_h2_s1_chipselect),            //                                .chipselect
		.REG_LED_s1_address                    (mm_interconnect_0_reg_led_s1_address),              //                      REG_LED_s1.address
		.REG_LED_s1_write                      (mm_interconnect_0_reg_led_s1_write),                //                                .write
		.REG_LED_s1_readdata                   (mm_interconnect_0_reg_led_s1_readdata),             //                                .readdata
		.REG_LED_s1_writedata                  (mm_interconnect_0_reg_led_s1_writedata),            //                                .writedata
		.REG_LED_s1_chipselect                 (mm_interconnect_0_reg_led_s1_chipselect),           //                                .chipselect
		.REG_M1_s1_address                     (mm_interconnect_0_reg_m1_s1_address),               //                       REG_M1_s1.address
		.REG_M1_s1_write                       (mm_interconnect_0_reg_m1_s1_write),                 //                                .write
		.REG_M1_s1_readdata                    (mm_interconnect_0_reg_m1_s1_readdata),              //                                .readdata
		.REG_M1_s1_writedata                   (mm_interconnect_0_reg_m1_s1_writedata),             //                                .writedata
		.REG_M1_s1_chipselect                  (mm_interconnect_0_reg_m1_s1_chipselect),            //                                .chipselect
		.REG_M2_s1_address                     (mm_interconnect_0_reg_m2_s1_address),               //                       REG_M2_s1.address
		.REG_M2_s1_write                       (mm_interconnect_0_reg_m2_s1_write),                 //                                .write
		.REG_M2_s1_readdata                    (mm_interconnect_0_reg_m2_s1_readdata),              //                                .readdata
		.REG_M2_s1_writedata                   (mm_interconnect_0_reg_m2_s1_writedata),             //                                .writedata
		.REG_M2_s1_chipselect                  (mm_interconnect_0_reg_m2_s1_chipselect),            //                                .chipselect
		.REG_S1_s1_address                     (mm_interconnect_0_reg_s1_s1_address),               //                       REG_S1_s1.address
		.REG_S1_s1_write                       (mm_interconnect_0_reg_s1_s1_write),                 //                                .write
		.REG_S1_s1_readdata                    (mm_interconnect_0_reg_s1_s1_readdata),              //                                .readdata
		.REG_S1_s1_writedata                   (mm_interconnect_0_reg_s1_s1_writedata),             //                                .writedata
		.REG_S1_s1_chipselect                  (mm_interconnect_0_reg_s1_s1_chipselect),            //                                .chipselect
		.REG_S2_s1_address                     (mm_interconnect_0_reg_s2_s1_address),               //                       REG_S2_s1.address
		.REG_S2_s1_write                       (mm_interconnect_0_reg_s2_s1_write),                 //                                .write
		.REG_S2_s1_readdata                    (mm_interconnect_0_reg_s2_s1_readdata),              //                                .readdata
		.REG_S2_s1_writedata                   (mm_interconnect_0_reg_s2_s1_writedata),             //                                .writedata
		.REG_S2_s1_chipselect                  (mm_interconnect_0_reg_s2_s1_chipselect),            //                                .chipselect
		.TIMER_s1_address                      (mm_interconnect_0_timer_s1_address),                //                        TIMER_s1.address
		.TIMER_s1_write                        (mm_interconnect_0_timer_s1_write),                  //                                .write
		.TIMER_s1_readdata                     (mm_interconnect_0_timer_s1_readdata),               //                                .readdata
		.TIMER_s1_writedata                    (mm_interconnect_0_timer_s1_writedata),              //                                .writedata
		.TIMER_s1_chipselect                   (mm_interconnect_0_timer_s1_chipselect),             //                                .chipselect
		.UART_s1_address                       (mm_interconnect_0_uart_s1_address),                 //                         UART_s1.address
		.UART_s1_write                         (mm_interconnect_0_uart_s1_write),                   //                                .write
		.UART_s1_read                          (mm_interconnect_0_uart_s1_read),                    //                                .read
		.UART_s1_readdata                      (mm_interconnect_0_uart_s1_readdata),                //                                .readdata
		.UART_s1_writedata                     (mm_interconnect_0_uart_s1_writedata),               //                                .writedata
		.UART_s1_begintransfer                 (mm_interconnect_0_uart_s1_begintransfer),           //                                .begintransfer
		.UART_s1_chipselect                    (mm_interconnect_0_uart_s1_chipselect)               //                                .chipselect
	);

	clock_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
