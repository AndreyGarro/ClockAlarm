// clock_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module clock_tb (
	);

	wire        clock_inst_clk_bfm_clk_clk;                     // clock_inst_clk_bfm:clk -> [clock_inst:clk_clk, clock_inst_reset_bfm:clk, clock_inst_timer_irq_bfm:clk, irq_mapper:clk]
	wire  [7:0] clock_inst_reg_h1_external_connection_export;   // clock_inst:reg_h1_external_connection_export -> clock_inst_reg_h1_external_connection_bfm:sig_export
	wire  [7:0] clock_inst_reg_h2_external_connection_1_export; // clock_inst:reg_h2_external_connection_1_export -> clock_inst_reg_h2_external_connection_1_bfm:sig_export
	wire  [7:0] clock_inst_reg_m1_external_connection_export;   // clock_inst:reg_m1_external_connection_export -> clock_inst_reg_m1_external_connection_bfm:sig_export
	wire  [7:0] clock_inst_reg_m2_external_connection_export;   // clock_inst:reg_m2_external_connection_export -> clock_inst_reg_m2_external_connection_bfm:sig_export
	wire  [7:0] clock_inst_reg_s1_external_connection_export;   // clock_inst:reg_s1_external_connection_export -> clock_inst_reg_s1_external_connection_bfm:sig_export
	wire  [7:0] clock_inst_reg_s2_external_connection_export;   // clock_inst:reg_s2_external_connection_export -> clock_inst_reg_s2_external_connection_bfm:sig_export
	wire        clock_inst_reset_bfm_reset_reset;               // clock_inst_reset_bfm:reset -> [clock_inst:reset_reset_n, clock_inst_timer_irq_bfm:reset, irq_mapper:reset]
	wire        irq_mapper_receiver0_irq;                       // clock_inst:timer_irq_irq -> irq_mapper:receiver0_irq
	wire  [0:0] clock_inst_timer_irq_bfm_irq_irq;               // irq_mapper:sender_irq -> clock_inst_timer_irq_bfm:irq

	clock clock_inst (
		.clk_clk                             (clock_inst_clk_bfm_clk_clk),                     //                          clk.clk
		.reg_h1_external_connection_export   (clock_inst_reg_h1_external_connection_export),   //   reg_h1_external_connection.export
		.reg_h2_external_connection_1_export (clock_inst_reg_h2_external_connection_1_export), // reg_h2_external_connection_1.export
		.reg_m1_external_connection_export   (clock_inst_reg_m1_external_connection_export),   //   reg_m1_external_connection.export
		.reg_m2_external_connection_export   (clock_inst_reg_m2_external_connection_export),   //   reg_m2_external_connection.export
		.reg_s1_external_connection_export   (clock_inst_reg_s1_external_connection_export),   //   reg_s1_external_connection.export
		.reg_s2_external_connection_export   (clock_inst_reg_s2_external_connection_export),   //   reg_s2_external_connection.export
		.reset_reset_n                       (clock_inst_reset_bfm_reset_reset),               //                        reset.reset_n
		.timer_irq_irq                       (irq_mapper_receiver0_irq)                        //                    timer_irq.irq
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) clock_inst_clk_bfm (
		.clk (clock_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm clock_inst_reg_h1_external_connection_bfm (
		.sig_export (clock_inst_reg_h1_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm clock_inst_reg_h2_external_connection_1_bfm (
		.sig_export (clock_inst_reg_h2_external_connection_1_export)  // conduit.export
	);

	altera_conduit_bfm clock_inst_reg_m1_external_connection_bfm (
		.sig_export (clock_inst_reg_m1_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm clock_inst_reg_m2_external_connection_bfm (
		.sig_export (clock_inst_reg_m2_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm clock_inst_reg_s1_external_connection_bfm (
		.sig_export (clock_inst_reg_s1_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm clock_inst_reg_s2_external_connection_bfm (
		.sig_export (clock_inst_reg_s2_external_connection_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) clock_inst_reset_bfm (
		.reset (clock_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (clock_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_avalon_interrupt_sink #(
		.ASSERT_HIGH_IRQ        (1),
		.AV_IRQ_W               (1),
		.ASYNCHRONOUS_INTERRUPT (0),
		.VHDL_ID                (0)
	) clock_inst_timer_irq_bfm (
		.clk   (clock_inst_clk_bfm_clk_clk),        //       clock_reset.clk
		.reset (~clock_inst_reset_bfm_reset_reset), // clock_reset_reset.reset
		.irq   (clock_inst_timer_irq_bfm_irq_irq)   //               irq.irq
	);

	altera_irq_mapper irq_mapper (
		.clk           (clock_inst_clk_bfm_clk_clk),        //       clk.clk
		.reset         (~clock_inst_reset_bfm_reset_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),          // receiver0.irq
		.sender_irq    (clock_inst_timer_irq_bfm_irq_irq)   //    sender.irq
	);

endmodule
